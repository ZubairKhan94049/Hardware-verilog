library verilog;
use verilog.vl_types.all;
entity buffer_stim is
end buffer_stim;
