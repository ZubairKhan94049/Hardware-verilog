library verilog;
use verilog.vl_types.all;
entity orgateusingnand_stim is
end orgateusingnand_stim;
