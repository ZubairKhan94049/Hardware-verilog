library verilog;
use verilog.vl_types.all;
entity \buffer\ is
    port(
        x               : in     vl_logic;
        y               : out    vl_logic
    );
end \buffer\;
